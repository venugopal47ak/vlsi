
module pg(input [3:0] d,output parity);
    assign parity=^d;
      endmodule
      
